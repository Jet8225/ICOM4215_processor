module decoder_4x16_neg(output reg [15:0] Y, input [3:0] X);
	always @(X)
		case(X)
			4'h0:	Y = 16'b1111111111111110;
			4'h1:	Y = 16'b1111111111111101;
			4'h2: 	Y = 16'b1111111111111011;
			4'h3:	Y = 16'b1111111111110111;
			4'h4:	Y = 16'b1111111111101111;
			4'h5:	Y = 16'b1111111111011111;
			4'h6: 	Y = 16'b1111111110111111;
			4'h7:	Y = 16'b1111111101111111;
			4'h8:	Y = 16'b1111111011111111;
			4'h9:	Y = 16'b1111110111111111;
			4'hA:	Y = 16'b1111101111111111;
			4'hB:	Y = 16'b1111011111111111;
			4'hC:	Y = 16'b1110111111111111;
			4'hD:	Y = 16'b1101111111111111;
			4'hE:	Y = 16'b1011111111111111;
			4'hF:	Y = 16'b0111111111111111;
		endcase
endmodule
